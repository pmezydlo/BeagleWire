module gpio (inout  [GPIO_WIDTH-1:0] io,
             input  [GPIO_WIDTH-1:0] dir,
             input  [GPIO_WIDTH-1:0] set,
             output [GPIO_WIDTH-1:0] get,

parameter GPIO_WIDTH = 32;

assign 

endmodule
